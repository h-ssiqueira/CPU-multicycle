LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY ULAExt IS
	PORT( ALUSrcA1,clock1		:IN	STD_LOGIC;
			ALUop1,ALUSrcB1	:IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
			A1, B1,PC1,Imed1 :IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
			ALUout1 		    :OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ULAExt;


ARCHITECTURE options OF ULAExt IS
COMPONENT ULA
PORT(
    ALUSrcA,clock		:IN	STD_LOGIC;
    ALUop,ALUSrcB	:IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
    A, B,PC,Imed	:IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
    ALUout 			:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;
BEGIN
    LUA: ULA PORT MAP (ALUSrcA1, clock1, ALUop1, ALUSrcB1, A1,B1, PC1,Imed1, ALUout1);
END options;
