LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PCATT IS
	PORT( PCWrite1,CLOCK1		:IN STD_LOGIC;
			ADDRESS		:IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
			ADDRESSATT	:BUFFER STD_LOGIC_VECTOR(7 DOWNTO 0));
END PCATT;

ARCHITECTURE options OF PCATT IS
BEGIN
	PROCESS(PCWrite1, ADDRESS,CLOCK1)
	BEGIN
	IF CLOCK1'EVENT AND CLOCK1 = '0' THEN
		 IF (PCWrite1 = '1' AND ADDRESS = "01000000") THEN
			ADDRESSATT <= "00000000";
		 ELSIF PCWrite1 = '1' THEN
			ADDRESSATT <= ADDRESS;
		END IF;
	END IF;
	END PROCESS;
END options;